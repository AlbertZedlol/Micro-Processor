//Instruction Memory
module InstructionMemory(
	input      [32 -1:0] Address, 
	
	output reg [32 -1:0] Instruction
);
	//maximum number of instructions: 2^{9-2+1}==256
	always @(*)
		case (Address[9:2])//Address[9:2] represents at most 256=2^{9-2+1}) instructions recorded in byte address, since address[1:0]are always zeros.(byte address)
			//Hexadecimal Machine Codes of Dijkstra Algorithm
			//codes generated with MARS compiler and python file process.py
          8'd0:	Instruction<=32'h24100000;
8'd1:	Instruction<=32'h3c014000;
8'd2:	Instruction<=32'h34310010;
8'd3:	Instruction<=32'h24120010;
8'd4:	Instruction<=32'h24080001;
8'd5:	Instruction<=32'h20050022;
8'd6:	Instruction<=32'h00054821;
8'd7:	Instruction<=32'h312a000f;
8'd8:	Instruction<=32'h000a5080;
8'd9:	Instruction<=32'h01505820;
8'd10:	Instruction<=32'h8d6c0000;
8'd11:	Instruction<=32'h00086a00;
8'd12:	Instruction<=32'h01ac7020;
8'd13:	Instruction<=32'hae2e0000;
8'd14:	Instruction<=32'h00094902;
8'd15:	Instruction<=32'h00084040;
8'd16:	Instruction<=32'h1512fff6;
8'd17:	Instruction<=32'h0000e021;
8'd18:	Instruction<=32'h0000e021;
8'd19:	Instruction<=32'h0000e021;
8'd20:	Instruction<=32'h0000e021;
8'd21:	Instruction<=32'h24080001;
8'd22:	Instruction<=32'h00054821;
8'd23:	Instruction<=32'h08000007;
8'd24:	Instruction<=32'h0000e021;
8'd25:	Instruction<=32'h0000e021;
8'd26:	Instruction<=32'h20080040;
8'd27:	Instruction<=32'h00082020;
8'd28:	Instruction<=32'h8d100000;
8'd29:	Instruction<=32'h21050004;
8'd30:	Instruction<=32'h0c000034;
8'd31:	Instruction<=32'h0000e021;
8'd32:	Instruction<=32'h0000e021;
8'd33:	Instruction<=32'h24080001;
8'd34:	Instruction<=32'h24080001;
8'd35:	Instruction<=32'h20090144;
8'd36:	Instruction<=32'h24050000;
8'd37:	Instruction<=32'h21290004;
8'd38:	Instruction<=32'h8d2a0000;
8'd39:	Instruction<=32'h00aa2820;
8'd40:	Instruction<=32'h21080001;
8'd41:	Instruction<=32'h0110082a;
8'd42:	Instruction<=32'h1420fffa;
8'd43:	Instruction<=32'h0000e021;
8'd44:	Instruction<=32'h0000e021;
8'd45:	Instruction<=32'h0000e021;
8'd46:	Instruction<=32'h0000e021;
8'd47:	Instruction<=32'h01004020;
8'd48:	Instruction<=32'h00084020;
8'd49:	Instruction<=32'h08000000;
8'd50:	Instruction<=32'h0000e021;
8'd51:	Instruction<=32'h0000e021;
8'd52:	Instruction<=32'h0000b021;
8'd53:	Instruction<=32'h22d60001;
8'd54:	Instruction<=32'h20010001;
8'd55:	Instruction<=32'h0001b822;
8'd56:	Instruction<=32'h20110144;
8'd57:	Instruction<=32'h00059021;
8'd58:	Instruction<=32'h20130194;
8'd59:	Instruction<=32'hae200000;
8'd60:	Instruction<=32'hae760000;
8'd61:	Instruction<=32'h00059021;
8'd62:	Instruction<=32'h00167821;
8'd63:	Instruction<=32'h01f0082a;
8'd64:	Instruction<=32'h10200011;
8'd65:	Instruction<=32'h0000e021;
8'd66:	Instruction<=32'h0000e021;
8'd67:	Instruction<=32'h0000e021;
8'd68:	Instruction<=32'h0000e021;
8'd69:	Instruction<=32'h000f6880;
8'd70:	Instruction<=32'h024d6820;
8'd71:	Instruction<=32'h8dad0000;
8'd72:	Instruction<=32'h000f4080;
8'd73:	Instruction<=32'h02284020;
8'd74:	Instruction<=32'had0d0000;
8'd75:	Instruction<=32'h000f5080;
8'd76:	Instruction<=32'h026a5020;
8'd77:	Instruction<=32'had400000;
8'd78:	Instruction<=32'h21ef0001;
8'd79:	Instruction<=32'h0800003f;
8'd80:	Instruction<=32'h0000e021;
8'd81:	Instruction<=32'h0000e021;
8'd82:	Instruction<=32'h00167821;
8'd83:	Instruction<=32'h01f0082a;
8'd84:	Instruction<=32'h1020006d;
8'd85:	Instruction<=32'h0000e021;
8'd86:	Instruction<=32'h0000e021;
8'd87:	Instruction<=32'h0000e021;
8'd88:	Instruction<=32'h0000e021;
8'd89:	Instruction<=32'h0017c021;
8'd90:	Instruction<=32'h00177021;
8'd91:	Instruction<=32'h0016c821;
8'd92:	Instruction<=32'h0330082a;
8'd93:	Instruction<=32'h10200028;
8'd94:	Instruction<=32'h0000e021;
8'd95:	Instruction<=32'h0000e021;
8'd96:	Instruction<=32'h0000e021;
8'd97:	Instruction<=32'h0000e021;
8'd98:	Instruction<=32'h00195080;
8'd99:	Instruction<=32'h026a5020;
8'd100:	Instruction<=32'h8d4c0000;
8'd101:	Instruction<=32'h00194880;
8'd102:	Instruction<=32'h02294820;
8'd103:	Instruction<=32'h8d2b0000;
8'd104:	Instruction<=32'h15800019;
8'd105:	Instruction<=32'h0000e021;
8'd106:	Instruction<=32'h0000e021;
8'd107:	Instruction<=32'h0000e021;
8'd108:	Instruction<=32'h0000e021;
8'd109:	Instruction<=32'h11770014;
8'd110:	Instruction<=32'h0000e021;
8'd111:	Instruction<=32'h0000e021;
8'd112:	Instruction<=32'h0000e021;
8'd113:	Instruction<=32'h0000e021;
8'd114:	Instruction<=32'h11d7000d;
8'd115:	Instruction<=32'h0000e021;
8'd116:	Instruction<=32'h0000e021;
8'd117:	Instruction<=32'h0000e021;
8'd118:	Instruction<=32'h0000e021;
8'd119:	Instruction<=32'h016e082a;
8'd120:	Instruction<=32'h14200007;
8'd121:	Instruction<=32'h0000e021;
8'd122:	Instruction<=32'h0000e021;
8'd123:	Instruction<=32'h0000e021;
8'd124:	Instruction<=32'h0000e021;
8'd125:	Instruction<=32'h08000082;
8'd126:	Instruction<=32'h0000e021;
8'd127:	Instruction<=32'h0000e021;
8'd128:	Instruction<=32'h000b7021;
8'd129:	Instruction<=32'h0019c021;
8'd130:	Instruction<=32'h23390001;
8'd131:	Instruction<=32'h0800005c;
8'd132:	Instruction<=32'h0000e021;
8'd133:	Instruction<=32'h0000e021;
8'd134:	Instruction<=32'h11d7003b;
8'd135:	Instruction<=32'h0000e021;
8'd136:	Instruction<=32'h0000e021;
8'd137:	Instruction<=32'h0000e021;
8'd138:	Instruction<=32'h0000e021;
8'd139:	Instruction<=32'h00185080;
8'd140:	Instruction<=32'h026a5020;
8'd141:	Instruction<=32'had560000;
8'd142:	Instruction<=32'h0016c821;
8'd143:	Instruction<=32'h0330082a;
8'd144:	Instruction<=32'h1020002d;
8'd145:	Instruction<=32'h0000e021;
8'd146:	Instruction<=32'h0000e021;
8'd147:	Instruction<=32'h0000e021;
8'd148:	Instruction<=32'h0000e021;
8'd149:	Instruction<=32'h00195080;
8'd150:	Instruction<=32'h026a5020;
8'd151:	Instruction<=32'h8d4c0000;
8'd152:	Instruction<=32'h001828c0;
8'd153:	Instruction<=32'h00b92820;
8'd154:	Instruction<=32'h00052880;
8'd155:	Instruction<=32'h0245e020;
8'd156:	Instruction<=32'h8f860000;
8'd157:	Instruction<=32'h1580001c;
8'd158:	Instruction<=32'h0000e021;
8'd159:	Instruction<=32'h0000e021;
8'd160:	Instruction<=32'h0000e021;
8'd161:	Instruction<=32'h0000e021;
8'd162:	Instruction<=32'h10d70017;
8'd163:	Instruction<=32'h0000e021;
8'd164:	Instruction<=32'h0000e021;
8'd165:	Instruction<=32'h0000e021;
8'd166:	Instruction<=32'h0000e021;
8'd167:	Instruction<=32'h00194880;
8'd168:	Instruction<=32'h02294820;
8'd169:	Instruction<=32'h8d240000;
8'd170:	Instruction<=32'h01c63820;
8'd171:	Instruction<=32'h1097000d;
8'd172:	Instruction<=32'h0000e021;
8'd173:	Instruction<=32'h0000e021;
8'd174:	Instruction<=32'h0000e021;
8'd175:	Instruction<=32'h0000e021;
8'd176:	Instruction<=32'h00e4082a;
8'd177:	Instruction<=32'h14200007;
8'd178:	Instruction<=32'h0000e021;
8'd179:	Instruction<=32'h0000e021;
8'd180:	Instruction<=32'h0000e021;
8'd181:	Instruction<=32'h0000e021;
8'd182:	Instruction<=32'h080000ba;
8'd183:	Instruction<=32'h0000e021;
8'd184:	Instruction<=32'h0000e021;
8'd185:	Instruction<=32'had270000;
8'd186:	Instruction<=32'h23390001;
8'd187:	Instruction<=32'h0800008f;
8'd188:	Instruction<=32'h0000e021;
8'd189:	Instruction<=32'h0000e021;
8'd190:	Instruction<=32'h21ef0001;
8'd191:	Instruction<=32'h08000053;
8'd192:	Instruction<=32'h0000e021;
8'd193:	Instruction<=32'h0000e021;
8'd194:	Instruction<=32'h03e00008;
8'd195:	Instruction<=32'h0000e021;
8'd196:	Instruction<=32'h0000e021;





            
            // 8'd0:	Instruction<=32'h08000001;
            // 8'd1:    Instruction<=32'h20080040;
            // 8'd2:    Instruction<=32'h00082020;
            // 8'd3:    Instruction<=32'h8d100000;
            // 8'd4:    Instruction<=32'h21050004;
            // 8'd5:    Instruction<=32'h0c000015;
            // 8'd6:    Instruction<=32'h24080001;
            // 8'd7:    Instruction<=32'h24080001;
            // 8'd8:    Instruction<=32'h20090144;
            // 8'd9:    Instruction<=32'h24050000;
            // 8'd10:    Instruction<=32'h21290004;
            // 8'd11:    Instruction<=32'h8d2a0000;
            // 8'd12:    Instruction<=32'h00aa2820;
            // 8'd13:    Instruction<=32'h21080001;
            // 8'd14:    Instruction<=32'h0110082a;
            // 8'd15:    Instruction<=32'h1420fffa;
            // 8'd16:    Instruction<=32'h01004020;
            // 8'd17:    Instruction<=32'h00084020;
            // 8'd18:    Instruction<=32'h24040000;
            // 8'd19:    Instruction<=32'h24020011;
            // 8'd20:    Instruction<=32'h0000000c;
            // 8'd21:    Instruction<=32'h0000b021;
            // 8'd22:    Instruction<=32'h22d60001;
            // 8'd23:    Instruction<=32'h20010001;
            // 8'd24:    Instruction<=32'h0001b822;
            // 8'd25:    Instruction<=32'h20110144;
            // 8'd26:    Instruction<=32'h00059021;
            // 8'd27:    Instruction<=32'h20130194;
            // 8'd28:    Instruction<=32'hae200000;
            // 8'd29:    Instruction<=32'hae760000;
            // 8'd30:    Instruction<=32'h00059021;
            // 8'd31:    Instruction<=32'h00167821;
            // 8'd32:    Instruction<=32'h01f0082a;
            // 8'd33:    Instruction<=32'h1020000b;
            // 8'd34:    Instruction<=32'h000f6880;
            // 8'd35:    Instruction<=32'h024d6820;
            // 8'd36:    Instruction<=32'h8dad0000;
            // 8'd37:    Instruction<=32'h000f4080;
            // 8'd38:    Instruction<=32'h02284020;
            // 8'd39:    Instruction<=32'had0d0000;
            // 8'd40:    Instruction<=32'h000f5080;
            // 8'd41:    Instruction<=32'h026a5020;
            // 8'd42:    Instruction<=32'had400000;
            // 8'd43:    Instruction<=32'h21ef0001;
            // 8'd44:    Instruction<=32'h08000020;
            // 8'd45:    Instruction<=32'h00167821;
            // 8'd46:    Instruction<=32'h01f0082a;
            // 8'd47:    Instruction<=32'h10200033;
            // 8'd48:    Instruction<=32'h0017c021;
            // 8'd49:    Instruction<=32'h00177021;
            // 8'd50:    Instruction<=32'h0016c821;
            // 8'd51:    Instruction<=32'h0330082a;
            // 8'd52:    Instruction<=32'h10200010;
            // 8'd53:    Instruction<=32'h00195080;
            // 8'd54:    Instruction<=32'h026a5020;
            // 8'd55:    Instruction<=32'h8d4c0000;
            // 8'd56:    Instruction<=32'h00194880;
            // 8'd57:    Instruction<=32'h02294820;
            // 8'd58:    Instruction<=32'h8d2b0000;
            // 8'd59:    Instruction<=32'h15800007;
            // 8'd60:    Instruction<=32'h11770006;
            // 8'd61:    Instruction<=32'h11d70003;
            // 8'd62:    Instruction<=32'h016e082a;
            // 8'd63:    Instruction<=32'h14200001;
            // 8'd64:    Instruction<=32'h08000043;
            // 8'd65:    Instruction<=32'h000b7021;
            // 8'd66:    Instruction<=32'h0019c021;
            // 8'd67:    Instruction<=32'h23390001;
            // 8'd68:    Instruction<=32'h08000033;
            // 8'd69:    Instruction<=32'h11d7001d;
            // 8'd70:    Instruction<=32'h00185080;
            // 8'd71:    Instruction<=32'h026a5020;
            // 8'd72:    Instruction<=32'had560000;
            // 8'd73:    Instruction<=32'h0016c821;
            // 8'd74:    Instruction<=32'h0330082a;
            // 8'd75:    Instruction<=32'h10200015;
            // 8'd76:    Instruction<=32'h00195080;
            // 8'd77:    Instruction<=32'h026a5020;
            // 8'd78:    Instruction<=32'h8d4c0000;
            // 8'd79:    Instruction<=32'h001828c0;
            // 8'd80:    Instruction<=32'h00b92820;
            // 8'd81:    Instruction<=32'h00052880;
            // 8'd82:    Instruction<=32'h0245e020;
            // 8'd83:    Instruction<=32'h8f860000;
            // 8'd84:    Instruction<=32'h1580000a;
            // 8'd85:    Instruction<=32'h10d70009;
            // 8'd86:    Instruction<=32'h00194880;
            // 8'd87:    Instruction<=32'h02294820;
            // 8'd88:    Instruction<=32'h8d240000;
            // 8'd89:    Instruction<=32'h01c63820;
            // 8'd90:    Instruction<=32'h10970003;
            // 8'd91:    Instruction<=32'h00e4082a;
            // 8'd92:    Instruction<=32'h14200001;
            // 8'd93:    Instruction<=32'h0800005f;
            // 8'd94:    Instruction<=32'had270000;
            // 8'd95:    Instruction<=32'h23390001;
            // 8'd96:    Instruction<=32'h0800004a;
            // 8'd97:    Instruction<=32'h21ef0001;
            // 8'd98:    Instruction<=32'h0800002e;
            // 8'd99:    Instruction<=32'h03e00008;
            default: Instruction <= 32'h00000000;
		endcase
		
endmodule
